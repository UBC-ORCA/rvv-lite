package opcodes;
  /////////////////////////////////////////////////////////////////////////////////
  //                                TEMPLATES                                    //
  /////////////////////////////////////////////////////////////////////////////////
  localparam [31:0] VALU_CFG        = 32'b?????????????????_???_?????_1010111;
  localparam [31:0] VALU_OPIVV      = 32'b??????_?_?????_?????_000_?????_1010111;
  localparam [31:0] VALU_OPFVV      = 32'b??????_?_?????_?????_001_?????_1010111;
  localparam [31:0] VALU_OPMVV      = 32'b??????_?_?????_?????_010_?????_1010111;
  localparam [31:0] VALU_OPIVI      = 32'b??????_?_?????_?????_011_?????_1010111;
  localparam [31:0] VALU_OPIVX      = 32'b??????_?_?????_?????_100_?????_1010111;
  localparam [31:0] VALU_OPFVF      = 32'b??????_?_?????_?????_101_?????_1010111;
  localparam [31:0] VALU_OPMVX      = 32'b??????_?_?????_?????_110_?????_1010111;
  localparam [31:0] VCFG            = 32'b?????????????????_111_?????_1010111;
  localparam [31:0] VLOAD           = 32'b???_?_??_?_?????_?????_???_?????_0000111;
  localparam [31:0] VSTORE          = 32'b???_?_??_?_?????_?????_???_?????_0100111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A1                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //a) vsetvli rd,rs1,vtypei # rd=VL=f(AVL), AVL=rs1, new vtype 
  //a) vsetivli rd,uimm,vtypei # rd=VL=f(AVL), AVL=uimm, new vtype 
  //a) vsetvl rd, rs1, rs2 # rd=VL=f(AVL), AVL=rs1, vtype=rs2 
  //a) vleEW.v vd,(rs1),vm # vector load, EEW=EW 
  //a) vseEW.v vs3,(rs1),vm # vector store, EEW=EW
  localparam [31:0] VSETVLI         = 32'b0????????????????_111_?????_1010111;
  localparam [31:0] VSETIVLI        = 32'b11???????????????_111_?????_1010111;
  localparam [31:0] VSETVL          = 32'b1000000??????????_111_?????_1010111;
  localparam [31:0] VLE_8_V         = 32'b???_0_00_?_00000_?????_000_?????_0000111;
  localparam [31:0] VLE_16_V        = 32'b???_0_00_?_00000_?????_101_?????_0000111;
  localparam [31:0] VLE_32_V        = 32'b???_0_00_?_00000_?????_110_?????_0000111;
  localparam [31:0] VLE_64_V        = 32'b???_0_00_?_00000_?????_111_?????_0000111;
  localparam [31:0] VSE_8_V         = 32'b???_0_00_?_00000_?????_000_?????_0100111;
  localparam [31:0] VSE_16_V        = 32'b???_0_00_?_00000_?????_101_?????_0100111;
  localparam [31:0] VSE_32_V        = 32'b???_0_00_?_00000_?????_110_?????_0100111;
  localparam [31:0] VSE_64_V        = 32'b???_0_00_?_00000_?????_111_?????_0100111;

  //b) vLOP.VXI vd,vs2,YY,vm # vd[i] = vs2[i] LOP YY 
  //b) vADDSUB.VXI vd,vs2,YY,vm # vd[i] = vs2[i] ADDSUB YY 
  //b) vrsub.XI vd,vs2,YY,vm # vd[i] = YY - vs2[i]
  //b) vid.v vd,vm # vd[i] = i 
  localparam [31:0] VAND_VV         = 32'b001001_?_?????_?????_000_?????_1010111;
  localparam [31:0] VAND_VX         = 32'b001001_?_?????_?????_100_?????_1010111;
  localparam [31:0] VAND_VI         = 32'b001001_?_?????_?????_011_?????_1010111;
  localparam [31:0] VOR_VV          = 32'b001010_?_?????_?????_000_?????_1010111;
  localparam [31:0] VOR_VX          = 32'b001010_?_?????_?????_100_?????_1010111;
  localparam [31:0] VOR_VI          = 32'b001010_?_?????_?????_011_?????_1010111;
  localparam [31:0] VXOR_VV         = 32'b001011_?_?????_?????_000_?????_1010111;
  localparam [31:0] VXOR_VX         = 32'b001011_?_?????_?????_100_?????_1010111;
  localparam [31:0] VXOR_VI         = 32'b001011_?_?????_?????_011_?????_1010111;
  localparam [31:0] VADD_VV         = 32'b000000_?_?????_?????_000_?????_1010111;
  localparam [31:0] VADD_VX         = 32'b000000_?_?????_?????_100_?????_1010111;
  localparam [31:0] VADD_VI         = 32'b000000_?_?????_?????_011_?????_1010111;
  localparam [31:0] VSUB_VV         = 32'b000010_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSUB_VX         = 32'b000010_?_?????_?????_100_?????_1010111;
  localparam [31:0] VRSUB_VX        = 32'b000011_?_?????_?????_100_?????_1010111;
  localparam [31:0] VRSUB_VI        = 32'b000011_?_?????_?????_011_?????_1010111;
  localparam [31:0] VID_V           = 32'b010100_?_00000_10001_010_?????_1010111;

  //c) vMINMAX{U}.VX vd,vs2,YY,vm # vd[i] = MINMAX{U}(vs2[i], YY) 
  localparam [31:0] VMINU_VV        = 32'b000100_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMINU_VX        = 32'b000100_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMIN_VV         = 32'b000101_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMIN_VX         = 32'b000101_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMAXU_VV        = 32'b000110_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMAXU_VX        = 32'b000110_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMAX_VV         = 32'b000111_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMAX_VX         = 32'b000111_?_?????_?????_100_?????_1010111;

  //d) vmMCMP.VXI vd,vs2,YY,vm # vd.m[i] = (vs2[i] MCMP YY) 
  //d) vmSLT.VX vd,vs2,YY,vm # vd.m[i] = (vs2[i] < YY) 
  //d) vmSGT.XI vd,vs2,YY,vm # vd.m[i] = (vs2[i] > YY) 
  //d) vmMOP.mm vd,vs2,vs1 # vd.m[i] = MOP(vs2.m[i],vs1.m[i])
  localparam [31:0] VMSEQ_VV        = 32'b011000_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSEQ_VX        = 32'b011000_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSEQ_VI        = 32'b011000_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMSNE_VV        = 32'b011001_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSNE_VX        = 32'b011001_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSNE_VI        = 32'b011001_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMSLE_VV        = 32'b011101_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSLE_VX        = 32'b011101_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSLE_VI        = 32'b011101_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMSLEU_VV       = 32'b011100_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSLEU_VX       = 32'b011100_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSLEU_VI       = 32'b011100_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMSLT_VV        = 32'b011011_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSLT_VX        = 32'b011011_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSGT_VX        = 32'b011111_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMSGT_VI        = 32'b011111_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMANDNOT_MM     = 32'b011000_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMAND_MM        = 32'b011001_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMOR_MM         = 32'b011010_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMXOR_MM        = 32'b011011_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMORNOT_MM      = 32'b011100_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMNAND_MM       = 32'b011101_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMNOR_MM        = 32'b011110_1_?????_?????_010_?????_1010111;
  localparam [31:0] VMXNOR_MM       = 32'b011111_1_?????_?????_010_?????_1010111;

  //e) vmv.v.VXI vd,YY # vd[i] = YY, XI modes: integer splat 
  //e) vmv.x.s rd,vs2 # x[rd] = vs2[0], scalar copy (vs1=0) 
  //e) vmv.s.x vd,rs1 # vd[0] = x[rs1], scalar copy (vs2=0) 
  localparam [31:0] VMV_VV          = 32'b010111_1_00000_?????_000_?????_1010111;
  localparam [31:0] VMV_VX          = 32'b010111_1_00000_?????_100_?????_1010111;
  localparam [31:0] VMV_VI          = 32'b010111_1_00000_?????_011_?????_1010111;
  localparam [31:0] VMV_SX          = 32'b010000_1_00000_?????_110_?????_1010111;
  localparam [31:0] VMV_XS          = 32'b010000_1_?????_00000_010_?????_1010111;

  //f) vmvKr.v vd,vs2 # whole-vec. reg. group copy EMUL=K 
  //f) vlKEW.v vd,(a0) # whole reg EMUL=K, VLEN/EW elements, ignores VL 
  //f) vsKr.v vd,(a1) # whole reg EMUL=K, VLEN bits, ignores VL
  localparam [31:0] VMV_1_R_V       = 32'b100111_1_?????_00000_011_?????_1010111;
  localparam [31:0] VMV_2_R_V       = 32'b100111_1_?????_00001_011_?????_1010111;
  localparam [31:0] VMV_4_R_V       = 32'b100111_1_?????_00011_011_?????_1010111;
  localparam [31:0] VMV_8_R_V       = 32'b100111_1_?????_00111_011_?????_1010111;
  localparam [31:0] VL_1_RE_8_V     = 32'b000_0_00_1_01000_?????_000_?????_0000111;
  localparam [31:0] VL_2_RE_16_V    = 32'b001_0_00_1_01000_?????_101_?????_0000111;
  localparam [31:0] VL_4_RE_32_V    = 32'b011_0_00_1_01000_?????_110_?????_0000111;
  localparam [31:0] VL_8_RE_64_V    = 32'b111_0_00_1_01000_?????_111_?????_0000111;
  localparam [31:0] VS_1_R_V        = 32'b000_0_00_1_01000_?????_000_?????_0100111;
  localparam [31:0] VS_2_R_V        = 32'b001_0_00_1_01000_?????_000_?????_0100111;
  localparam [31:0] VS_4_R_V        = 32'b011_0_00_1_01000_?????_000_?????_0100111;
  localparam [31:0] VS_8_R_V        = 32'b111_0_00_1_01000_?????_000_?????_0100111;

  //g) vslide1up.vx vd,vs2,rs1,vm # vd[i+1]=vs2[i], vd[0]=X[rs1] 
  //g) vslide1down.vx vd,vs2,rs1,vm # vd[i]=vs2[i+1], vd[L]=X[rs1]
  localparam [31:0] VSLIDE1UP_VX    = 32'b001110_?_?????_?????_110_?????_1010111;
  localparam [31:0] VSLIDE1DOWN_VX  = 32'b001111_?_?????_?????_110_?????_1010111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A2                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vwADDSUB{U}.VX vd,vs2,YY,vm # vd[i] = vs2[i] ADDSUB{U} YY
  localparam [31:0] VWADDU_VV       = 32'b110000_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWADDU_VX       = 32'b110000_?_?????_?????_110_?????_1010111;
  localparam [31:0] VWADD_VV        = 32'b110001_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWADD_VX        = 32'b110001_?_?????_?????_110_?????_1010111;
  localparam [31:0] VWSUBU_VV       = 32'b110010_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWSUBU_VX       = 32'b110010_?_?????_?????_110_?????_1010111;
  localparam [31:0] VWSUB_VV        = 32'b110011_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWSUB_VX        = 32'b110011_?_?????_?????_110_?????_1010111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A3                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vredROP.vs vd,vs2,vs1,vm # vd[0]=ROP(vs1[0],vs2[*])
  localparam [31:0] VREDSUM_VS      = 32'b000000_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDAND_VS      = 32'b000001_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDOR_VS       = 32'b000010_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDXOR_VS      = 32'b000011_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDMINU_VS     = 32'b000100_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDMIN_VS      = 32'b000101_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDMAXU_VS     = 32'b000110_?_?????_?????_010_?????_1010111;
  localparam [31:0] VREDMAX_VS      = 32'b000111_?_?????_?????_010_?????_1010111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A4                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //a) vmul.VX vd,vs2,YY,vm # vd[i] = LSB(vs2[i] * YY) (8/16/32b) 
  //a) vsll.VXI vd,vs2,ZZ,vm # vd[i] = vs2[i] << YY (8/16/32b) 
  localparam [31:0] VMUL_VV         = 32'b100101_?_?????_?????_010_?????_1010111;
  localparam [31:0] VMUL_VX         = 32'b100101_?_?????_?????_110_?????_1010111;
  localparam [31:0] VSLL_VV         = 32'b100101_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSLL_VX         = 32'b100101_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSLL_VI         = 32'b100101_?_?????_?????_011_?????_1010111;

  //b) vsr{l/a}.VXI vd,vs2,ZZ,vm # vd[i] = vs2[i] {>}>> YY (8/16b) 
  //b) vMULH.VX vd,vs2,YY,vm # vd[i] = MSB(vs2[i] * YY) (8/16b) 
  //c) vsr{l/a}.VXI vd,vs2,ZZ,vm # vd[i] = vs2[i] {>}>> YY (32b) 
  //c) vMULH.VX vd,vs2,YY,vm # vd[i] = MSB(vs2[i] * YY) (32b)
  localparam [31:0] VSRL_VV         = 32'b101000_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSRL_VX         = 32'b101000_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSRL_VI         = 32'b101000_?_?????_?????_011_?????_1010111;
  localparam [31:0] VSRA_VV         = 32'b101001_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSRA_VX         = 32'b101001_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSRA_VI         = 32'b101001_?_?????_?????_011_?????_1010111;
  localparam [31:0] VMULH_VV        = 32'b100111_?_?????_?????_010_?????_1010111;
  localparam [31:0] VMULH_VX        = 32'b100111_?_?????_?????_110_?????_1010111;

  //d) vwMUL.VX vd,vs2,YY,vm # vd[i] = vs2[i] * YY (8/16/32b) 
  //d) vwmulsu.VX vd,vs2,YY,vm # vd[i] = vs2[i] S*U YY (8/16/32b) 
  //d) vnsrl.wX vd,vs2,x0,vm # vd[i] = vs2[i] (16/32/64b)
  localparam [31:0] VWMUL_VV        = 32'b111011_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWMUL_VX        = 32'b111011_?_?????_?????_110_?????_1010111;
  localparam [31:0] VWMULSU_VV      = 32'b111010_?_?????_?????_010_?????_1010111;
  localparam [31:0] VWMULSU_VX      = 32'b111010_?_?????_?????_110_?????_1010111;
  localparam [31:0] VNSRL_VV        = 32'b101100_?_?????_?????_000_?????_1010111;
  localparam [31:0] VNSRL_VX        = 32'b101100_?_?????_?????_100_?????_1010111;
  localparam [31:0] VNSRL_VI        = 32'b101100_?_?????_?????_011_?????_1010111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A5                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vslideup.XI vd,vs2,ZZ,vm # vd[i+ZZ] = vs2[i] 
  //vslidedown.XI vd,vs2,ZZ,vm # vd[i] = vs2[i+ZZ]
  localparam [31:0] VSLIDEUP_VX     = 32'b001110_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSLIDEUP_VI     = 32'b001110_?_?????_?????_011_?????_1010111;
  localparam [31:0] VSLIDEDOWN_VX   = 32'b001111_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSLIDEDOWN_VI   = 32'b001111_?_?????_?????_011_?????_1010111;

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A6                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vmul.VX vd,vs2,YY,vm # vd[i] = LSB(vs2[i] * YY) 
  //vsll.VXI vd,vs2,ZZ,vm # vd[i] = vs2[i] << YY 
  //vsr{l/a}.VXI vd,vs2,ZZ,vm # vd[i] = vs2[i] {>}>> YY

  /* 64-bit multiplication and shifting instructions from A4 */

  /////////////////////////////////////////////////////////////////////////////////
  //                                    A7                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vaADDSUB{U}.VX vd, vs2, YY, vm # round_US(vs2[i] ADDSUB{U} YY, 1) 
  //vsmul.VX vd, vs2, YY, vm # vd[i]=clip(round_S(vs2[i]*YY,SEW-1)) (no 64b) 
  //vssr{l/a}.VXI vd, vs2, ZZ, vm # vd[i]=round_{U}S(vs2[i],ZZ)
  localparam [31:0] VAADDU_VV       = 32'b001000_?_?????_?????_010_?????_1010111;
  localparam [31:0] VAADDU_VX       = 32'b001000_?_?????_?????_110_?????_1010111;
  localparam [31:0] VAADD_VV        = 32'b001001_?_?????_?????_010_?????_1010111;
  localparam [31:0] VAADD_VX        = 32'b001001_?_?????_?????_110_?????_1010111;
  localparam [31:0] VASUBU_VV       = 32'b001010_?_?????_?????_010_?????_1010111;
  localparam [31:0] VASUBU_VX       = 32'b001010_?_?????_?????_110_?????_1010111;
  localparam [31:0] VASUB_VV        = 32'b001011_?_?????_?????_010_?????_1010111;
  localparam [31:0] VASUB_VX        = 32'b001011_?_?????_?????_110_?????_1010111;
  localparam [31:0] VSMUL_VV        = 32'b100111_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSMUL_VX        = 32'b100111_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSSRL_VV        = 32'b101010_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSSRL_VX        = 32'b101010_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSSRL_VI        = 32'b101010_?_?????_?????_011_?????_1010111;
  localparam [31:0] VSSRA_VV        = 32'b101011_?_?????_?????_000_?????_1010111;
  localparam [31:0] VSSRA_VX        = 32'b101011_?_?????_?????_100_?????_1010111;
  localparam [31:0] VSSRA_VI        = 32'b101011_?_?????_?????_011_?????_1010111;
  
  /////////////////////////////////////////////////////////////////////////////////
  //                                    B1                                       //
  /////////////////////////////////////////////////////////////////////////////////

  //vlm.v vd, (rs1) # ld mask of ceil(vl/8) bytes 
  //vsm.v vs3,(rs1) # st mask of ceil(vl/8) bytes 
  //vadc.VXIm vd,vs2,YY,v0 # vd[i]=vs2[i]+vs1[i]+v0.m[i] 
  //vmadc.VXm vd,vs2,YY,v0 # vd.m[i]=cout(vs2[i]+vs1[i]+v0.m[i]) 
  //vmadc.VXI vd,vs2,YY # vd.m[i]=cout(vs2[i]+vs1[i]) 
  //vsbc.VXm vd,vs2,YY,v0 # vd[i]=vs2[i]-vs1[i]-v0.m[i] 
  //vmsbc.VXm vd,vs2,YY,v0 # vd.m[i]=brrw(vs2[i]-vs1[i]-v0.m[i]) 
  //vmsbc.VX vd,vs2,YY # vd.m[i]=brrw(vs2[i]-vs1[i]) 
  //vcpop.m rd,vs2,vm # x[rd] = sum(vs2.m[i]), count bits 
  //vfirst.m rd,vs2,vm # x[rd] = idx_of_first_one(vs2.m) 
  //vmerge.VXIm vd,vs2,YY,v0 # vd[i] = v0.m[i] ? YY : vs2[i]
  localparam [31:0] VLM_V           = 32'b000_0_00_1_01011_?????_000_?????_0000111;
  localparam [31:0] VSM_V           = 32'b000_0_00_1_01011_?????_000_?????_0100111;
  localparam [31:0] VCPOP_M         = 32'b010000_?_?????_10000_010_?????_1010111;
  localparam [31:0] VFIRST_M        = 32'b010000_?_?????_10001_010_?????_1010111;
  localparam [31:0] VMERGE_VV       = 32'b010111_0_?????_?????_000_?????_1010111;
  localparam [31:0] VMERGE_VX       = 32'b010111_0_?????_?????_100_?????_1010111;
  localparam [31:0] VMERGE_VI       = 32'b010111_0_?????_?????_011_?????_1010111;
  localparam [31:0] VADC_VV         = 32'b010000_0_?????_?????_000_?????_1010111;
  localparam [31:0] VADC_VX         = 32'b010000_0_?????_?????_100_?????_1010111;
  localparam [31:0] VADC_VI         = 32'b010000_0_?????_?????_011_?????_1010111;
  localparam [31:0] VMADC_VV        = 32'b010001_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMADC_VX        = 32'b010001_?_?????_?????_100_?????_1010111;
  localparam [31:0] VMADC_VI        = 32'b010001_?_?????_?????_011_?????_1010111;
  localparam [31:0] VSBC_VV         = 32'b010010_0_?????_?????_000_?????_1010111;
  localparam [31:0] VSBC_VX         = 32'b010010_0_?????_?????_100_?????_1010111;
  localparam [31:0] VMSBC_VV        = 32'b010011_?_?????_?????_000_?????_1010111;
  localparam [31:0] VMSBC_VX        = 32'b010011_?_?????_?????_100_?????_1010111;

  typedef struct packed {
    logic [3-1:0] nf;
    logic mew;
    logic [2-1:0] mop;
    logic vm;
    logic [5-1:0] lumop;
    logic [5-1:0] rs1_addr;
    logic [3-1:0] width;
    logic [5-1:0] vd_addr;
    logic [7-1:0] opcode;
  } vload_instruction_t;

  typedef struct packed {
    logic [3-1:0] nf;
    logic mew;
    logic [2-1:0] mop;
    logic vm;
    logic [5-1:0] sumop;
    logic [5-1:0] rs1_addr;
    logic [3-1:0] width;
    logic [5-1:0] vs3_addr;
    logic [7-1:0] opcode;
  } vstore_instruction_t;

  typedef struct packed {
      logic [6-1:0] fn6;
      logic vm;
      logic [5-1:0] vs2_addr;
      logic [5-1:0] vs1_addr;
      logic [3-1:0] fn3;
      logic [5-1:0] vd_addr;
      logic [7-1:0] opcode;
  } valu_instruction_t;

  typedef struct packed {
    logic [7-1:0] fn7;
    logic [5-1:0] rs2_addr;
    logic [5-1:0] rs1_addr;
    logic [3-1:0] fn3;
    logic [5-1:0] rd_addr;
    logic [7-1:0] opcode;
  } vcfg_instruction_t;


  typedef struct packed {
    logic vill;
    logic [23-1:0] zeros;
    logic vma;
    logic vta;
    logic [3-1:0] vsew;
    logic [3-1:0] vlmul;
  } vtype_t;

endpackage
